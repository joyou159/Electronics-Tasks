
module posedge_detector(
    i_sig,
    i_clk,
    o_pe
);

    input i_sig;     // Input signal
    input i_clk;     // Clock signal

    output o_pe;     // Output signal indicating positive edge detection

    reg sig_delayed; // Internal register to store delayed input signal

    always @ (posedge i_clk) begin
        sig_delayed <= i_sig;  // Store the current input signal value on the positive edge of the clock
    end

    assign o_pe = i_sig & ~sig_delayed;  // Compare the current input signal with the delayed signal to detect positive edges

endmodule

/*In this code, posedge_detector is a module that detects positive edges on the i_sig input signal using the i_clk clock signal. 
Here are the explanations of the different sections and signals in the code:

input i_sig; and input i_clk; declare the input signals i_sig and i_clk.
output o_pe; declares the output signal o_pe, which indicates the detection of a positive edge.
reg sig_delayed; declares an internal register sig_delayed to store the delayed input signal value.
The always @ (posedge i_clk) block is sensitive to the positive edge of the clock signal i_clk.
Inside the always block, sig_delayed <= i_sig; assigns the current value of i_sig to sig_delayed on the positive edge of the clock.
assign o_pe = i_sig & ~sig_delayed; assigns the output o_pe the logical AND between the current i_sig and the negation of sig_delayed.
This results in a high output when a positive edge is detected.
This code captures the input signal value on the positive edge of the clock and compares it with the delayed value to determine positive edge detection.
The result is stored in the o_pe output signal.*/